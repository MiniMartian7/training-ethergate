package
    typedef enum bit [2:0] {WRITE = 'b101, READ = 'b110, IDLE = 'b100, ILLEGAL = 'b111, RESET = 'b000} e_operation;
endpackage