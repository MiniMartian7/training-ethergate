//  Interface: sif_i
//
interface sif_i #(
        <parameter_list>
    )(
        <port_list>
    );

    
endinterface: sif_i
