`include "sif_interface.sv"

module TB(sif_i tb_i);
    
endmodule : TB