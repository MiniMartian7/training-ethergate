module test (
    input logic [1:0] grant,
    output logic [1:0] request,
    output logic rst,
    input logic clk
);

initial begin
    @(posedge clk) request <= 2'b01;
    $display("@%0t: Drove req = 01", $time);
    repeat (2) @(posedge clk);
    if(grant != 2'b01) 
        $display("@%0t: a1: grant != 2'b01", $time);
    $finish;
end
endmodule