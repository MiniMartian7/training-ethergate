class enviroment;
    
endclass //enviroment