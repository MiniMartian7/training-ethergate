package
    typedef enum bit [2:0] {WRITE = 'b110, READ = 'b101, IDLE = 'b100, ILLEGAL = 'b111, RESET = 'b000} E_Operation;
endpackage