
class operation;
    logic [3:0] code;

    function new(logic [3:0] toDo);
      code = toDo;
    endfunction

    
endclass //operation

