module mem(
    clk_mem,
    rst_mem,
    
    en_in,
    digit_in,
    line_in,

    line_out
);

input clk_mem, rst_mem, en_in;
input [3:0] digit_in;

input [4:0] line_in;

output [31:0] line_out;

reg [31:0] line_out_d, line_out_ff;

reg [31:0] mem_nr_0 [0:31];
wire [31:0] buffer_0;

reg [31:0] mem_nr_1 [0:31];
wire [31:0] buffer_1;


reg [31:0] mem_nr_2 [0:31];
wire [31:0] buffer_2;


reg [31:0] mem_nr_3 [0:31];
wire [31:0] buffer_3; 


reg [31:0] mem_nr_4 [0:31]; 
wire [31:0] buffer_4;


reg [31:0] mem_nr_5 [0:31];
wire [31:0] buffer_5;


reg [31:0] mem_nr_6 [0:31];
wire [31:0] buffer_6;


reg [31:0] mem_nr_7 [0:31];
wire [31:0] buffer_7;


reg [31:0] mem_nr_8 [0:31];
wire [31:0] buffer_8;


reg [31:0] mem_nr_9 [0:31];
wire [31:0] buffer_9;


parameter ZERO = 'd0;
parameter ONE = 'd1;
parameter TWO = 'd2;
parameter THREE = 'd3;
parameter FOUR = 'd4;
parameter FIVE = 'd5;
parameter SIX = 'd6;
parameter SEVEN = 'd7;
parameter EIGTH = 'd8;
parameter NINE = 'd9;
parameter TEN = 'd10;

parameter NULL = 'b1111;

parameter ENABLE = 1;
parameter DISABLE = 0;
parameter RESET = 0;


always @(posedge clk_mem or posedge rst_mem) begin
    if(rst_mem) begin

        line_out_ff <= RESET;

        mem_nr_0[0] <= 32'b11111111111111111111111111111111;
        mem_nr_0[1] <= 32'b11111111111111111111111111111111;
        mem_nr_0[2] <= 32'b11111111111111111111111111111111;
        mem_nr_0[3] <= 32'b11111100000000000000000000111111;
        mem_nr_0[4] <= 32'b11111100000000000000000000111111;
        mem_nr_0[5] <= 32'b11111100000000000000000000111111;
        mem_nr_0[6] <= 32'b11111100000000000000000000111111;
        mem_nr_0[7] <= 32'b11111100000000000000000000111111;
        mem_nr_0[8] <= 32'b11111100000000000000000000111111;
        mem_nr_0[9] <= 32'b11111100000000000000000000111111;
        mem_nr_0[10] <= 32'b11111100000000000000000000111111;
        mem_nr_0[11] <= 32'b11111100000000000000000000111111;
        mem_nr_0[12] <= 32'b11111100000000000000000000111111;
        mem_nr_0[13] <= 32'b11111100000000000000000000111111;
        mem_nr_0[14] <= 32'b11111100000000000000000000111111;
        mem_nr_0[15] <= 32'b11111100000000000000000000111111;
        mem_nr_0[16] <= 32'b11111100000000000000000000111111;
        mem_nr_0[17] <= 32'b11111100000000000000000000111111;
        mem_nr_0[18] <= 32'b11111100000000000000000000111111;
        mem_nr_0[19] <= 32'b11111100000000000000000000111111;
        mem_nr_0[20] <= 32'b11111100000000000000000000111111;
        mem_nr_0[21] <= 32'b11111100000000000000000000111111;
        mem_nr_0[22] <= 32'b11111100000000000000000000111111;
        mem_nr_0[23] <= 32'b11111100000000000000000000111111;
        mem_nr_0[24] <= 32'b11111100000000000000000000111111;
        mem_nr_0[25] <= 32'b11111100000000000000000000111111;
        mem_nr_0[26] <= 32'b11111100000000000000000000111111;
        mem_nr_0[27] <= 32'b11111100000000000000000000111111;
        mem_nr_0[28] <= 32'b11111100000000000000000000111111;
        mem_nr_0[29] <= 32'b11111111111111111111111111111111;
        mem_nr_0[30] <= 32'b11111111111111111111111111111111;
        mem_nr_0[31] <= 32'b11111111111111111111111111111111;

mem_nr_1[0] = 32'b00000000000000000000000111111111;
mem_nr_1[1] = 32'b00000000000000000000011111111111;
mem_nr_1[2] = 32'b00000000000000000001111111111111;
mem_nr_1[3] = 32'b00000000000000000111111111111111;
mem_nr_1[4] = 32'b00000000000000011111111100111111;
mem_nr_1[5] = 32'b00000000000001111111110000111111;
mem_nr_1[6] = 32'b00000000000000000000000000111111;
mem_nr_1[7] = 32'b00000000000000000000000000111111;
mem_nr_1[8] = 32'b00000000000000000000000000111111;
mem_nr_1[9] = 32'b00000000000000000000000000111111;
mem_nr_1[10] = 32'b00000000000000000000000000111111;
mem_nr_1[11] = 32'b00000000000000000000000000111111;
mem_nr_1[12] = 32'b00000000000000000000000000111111;
mem_nr_1[13] = 32'b00000000000000000000000000111111;
mem_nr_1[14] = 32'b00000000000000000000000000111111;
mem_nr_1[15] = 32'b00000000000000000000000000111111;
mem_nr_1[16] = 32'b00000000000000000000000000111111;
mem_nr_1[17] = 32'b00000000000000000000000000111111;
mem_nr_1[18] = 32'b00000000000000000000000000111111;
mem_nr_1[19] = 32'b00000000000000000000000000111111;
mem_nr_1[20] = 32'b00000000000000000000000000111111;
mem_nr_1[21] = 32'b00000000000000000000000000111111;
mem_nr_1[22] = 32'b00000000000000000000000000111111;
mem_nr_1[23] = 32'b00000000000000000000000000111111;
mem_nr_1[24] = 32'b00000000000000000000000000111111;
mem_nr_1[25] = 32'b00000000000000000000000000111111;
mem_nr_1[26] = 32'b00000000000000000000000000111111;
mem_nr_1[27] = 32'b00000000000000000000000000111111;
mem_nr_1[28] = 32'b00000000000000000000000000111111;
mem_nr_1[29] = 32'b00000000000000000000000000111111;
mem_nr_1[30] = 32'b00000000000000000000000000111111;
mem_nr_1[31] = 32'b00000000000000000000000000111111;


mem_nr_2[0] <= 32'b11111111111111111111111111111111;
mem_nr_2[1] <= 32'b11111111111111111111111111111111;
mem_nr_2[2] <= 32'b11111111111111111111111111111111;
mem_nr_2[3] <= 32'b00000000000000000000000000111111;
mem_nr_2[4] <= 32'b00000000000000000000000000111111;
mem_nr_2[5] <= 32'b00000000000000000000000000111111;
mem_nr_2[6] <= 32'b00000000000000000000000000111111;
mem_nr_2[7] <= 32'b00000000000000000000000000111111;
mem_nr_2[8] <= 32'b00000000000000000000000000111111;
mem_nr_2[9] <= 32'b00000000000000000000000000111111;
mem_nr_2[10] <= 32'b00000000000000000000000000111111;
mem_nr_2[11] <= 32'b00000000000000000000000000111111;
mem_nr_2[12] <= 32'b00000000000000000000000000111111;
mem_nr_2[13] <= 32'b11111111111111111111111111111111;
mem_nr_2[14] <= 32'b11111111111111111111111111111111;
mem_nr_2[15] <= 32'b11111111111111111111111111111111;
mem_nr_2[16] <= 32'b11111111111111111111111111111111;
mem_nr_2[17] <= 32'b11111111111111111111111111111111;
mem_nr_2[18] <= 32'b11111100000000000000000000000000;
mem_nr_2[19] <= 32'b11111100000000000000000000000000;
mem_nr_2[20] <= 32'b11111100000000000000000000000000;
mem_nr_2[21] <= 32'b11111100000000000000000000000000;
mem_nr_2[22] <= 32'b11111100000000000000000000000000;
mem_nr_2[23] <= 32'b11111100000000000000000000000000;
mem_nr_2[24] <= 32'b11111100000000000000000000000000;
mem_nr_2[25] <= 32'b11111100000000000000000000000000;
mem_nr_2[26] <= 32'b11111100000000000000000000000000;
mem_nr_2[27] <= 32'b11111100000000000000000000000000;
mem_nr_2[28] <= 32'b11111100000000000000000000000000;
mem_nr_2[29] <= 32'b11111111111111111111111111111111;
mem_nr_2[30] <= 32'b11111111111111111111111111111111;
mem_nr_2[31] <= 32'b11111111111111111111111111111111;


mem_nr_3[0] <= 32'b11111111111111111111111111111111;
mem_nr_3[1] <= 32'b11111111111111111111111111111111;
mem_nr_3[2] <= 32'b11111111111111111111111111111111;
mem_nr_3[3] <= 32'b00000000000000000000000000111111;
mem_nr_3[4] <= 32'b00000000000000000000000000111111;
mem_nr_3[5] <= 32'b00000000000000000000000000111111;
mem_nr_3[6] <= 32'b00000000000000000000000000111111;
mem_nr_3[7] <= 32'b00000000000000000000000000111111;
mem_nr_3[8] <= 32'b00000000000000000000000000111111;
mem_nr_3[9] <= 32'b00000000000000000000000000111111;
mem_nr_3[10] <= 32'b00000000000000000000000000111111;
mem_nr_3[11] <= 32'b00000000000000000000000000111111;
mem_nr_3[12] <= 32'b00000000000000000000000000111111;
mem_nr_3[13] <= 32'b11111111111111111111111111111111;
mem_nr_3[14] <= 32'b11111111111111111111111111111111;
mem_nr_3[15] <= 32'b11111111111111111111111111111111;
mem_nr_3[16] <= 32'b11111111111111111111111111111111;
mem_nr_3[17] <= 32'b11111111111111111111111111111111;
mem_nr_3[18] <= 32'b00000000000000000000000000111111;
mem_nr_3[19] <= 32'b00000000000000000000000000111111;
mem_nr_3[20] <= 32'b00000000000000000000000000111111;
mem_nr_3[21] <= 32'b00000000000000000000000000111111;
mem_nr_3[22] <= 32'b00000000000000000000000000111111;
mem_nr_3[23] <= 32'b00000000000000000000000000111111;
mem_nr_3[24] <= 32'b00000000000000000000000000111111;
mem_nr_3[25] <= 32'b00000000000000000000000000111111;
mem_nr_3[26] <= 32'b00000000000000000000000000111111;
mem_nr_3[27] <= 32'b00000000000000000000000000111111;
mem_nr_3[28] <= 32'b00000000000000000000000000111111;
mem_nr_3[29] <= 32'b11111111111111111111111111111111;
mem_nr_3[30] <= 32'b11111111111111111111111111111111;
mem_nr_3[31] <= 32'b11111111111111111111111111111111;

mem_nr_4[0] <= 32'b11111100000000000000000000000000;
mem_nr_4[1] <= 32'b11111100000000000000000000000000;
mem_nr_4[2] <= 32'b11111100000000000000000000000000;
mem_nr_4[3] <= 32'b11111100000000000000000000000000;
mem_nr_4[4] <= 32'b11111100000000000000000000000000;
mem_nr_4[5] <= 32'b11111100000000000000000000000000;
mem_nr_4[6] <= 32'b11111100000000000000000000000000;
mem_nr_4[7] <= 32'b11111100000000000000000000000000;
mem_nr_4[8] <= 32'b11111100000000000000000000000000;
mem_nr_4[9] <= 32'b11111100000000000000000000000000;
mem_nr_4[10] <= 32'b11111100000000000000000000000000;
mem_nr_4[11] <= 32'b11111100000000000000000000000000;
mem_nr_4[12] <= 32'b11111100000000000000000000000000;
mem_nr_4[13] <= 32'b11111111111111111111111111111111;
mem_nr_4[14] <= 32'b11111111111111111111111111111111;
mem_nr_4[15] <= 32'b11111111111111111111111111111111;
mem_nr_4[16] <= 32'b11111111111111111111111111111111;
mem_nr_4[17] <= 32'b11111111111111111111111111111111;
mem_nr_4[18] <= 32'b00000000000000000000000000111111;
mem_nr_4[19] <= 32'b00000000000000000000000000111111;
mem_nr_4[20] <= 32'b00000000000000000000000000111111;
mem_nr_4[21] <= 32'b00000000000000000000000000111111;
mem_nr_4[22] <= 32'b00000000000000000000000000111111;
mem_nr_4[23] <= 32'b00000000000000000000000000111111;
mem_nr_4[24] <= 32'b00000000000000000000000000111111;
mem_nr_4[25] <= 32'b00000000000000000000000000111111;
mem_nr_4[26] <= 32'b00000000000000000000000000111111;
mem_nr_4[27] <= 32'b00000000000000000000000000111111;
mem_nr_4[28] <= 32'b00000000000000000000000000111111;
mem_nr_4[29] <= 32'b00000000000000000000000000111111;
mem_nr_4[30] <= 32'b00000000000000000000000000111111;
mem_nr_4[31] <= 32'b00000000000000000000000000111111;


mem_nr_5[0] <= 32'b11111111111111111111111111111111;
mem_nr_5[1] <= 32'b11111111111111111111111111111111;
mem_nr_5[2] <= 32'b11111111111111111111111111111111;
mem_nr_5[3] <= 32'b11111100000000000000000000000000;
mem_nr_5[4] <= 32'b11111100000000000000000000000000;
mem_nr_5[5] <= 32'b11111100000000000000000000000000;
mem_nr_5[6] <= 32'b11111100000000000000000000000000;
mem_nr_5[7] <= 32'b11111100000000000000000000000000;
mem_nr_5[8] <= 32'b11111100000000000000000000000000;
mem_nr_5[9] <= 32'b11111100000000000000000000000000;
mem_nr_5[10] <= 32'b11111100000000000000000000000000;
mem_nr_5[11] <= 32'b11111100000000000000000000000000;
mem_nr_5[12] <= 32'b11111100000000000000000000000000;
mem_nr_5[13] <= 32'b11111111111111111111111111111111;
mem_nr_5[14] <= 32'b11111111111111111111111111111111;
mem_nr_5[15] <= 32'b11111111111111111111111111111111;
mem_nr_5[16] <= 32'b11111111111111111111111111111111;
mem_nr_5[17] <= 32'b11111111111111111111111111111111;
mem_nr_5[18] <= 32'b00000000000000000000000000111111;
mem_nr_5[19] <= 32'b00000000000000000000000000111111;
mem_nr_5[20] <= 32'b00000000000000000000000000111111;
mem_nr_5[21] <= 32'b00000000000000000000000000111111;
mem_nr_5[22] <= 32'b00000000000000000000000000111111;
mem_nr_5[23] <= 32'b00000000000000000000000000111111;
mem_nr_5[24] <= 32'b00000000000000000000000000111111;
mem_nr_5[25] <= 32'b00000000000000000000000000111111;
mem_nr_5[26] <= 32'b00000000000000000000000000111111;
mem_nr_5[27] <= 32'b00000000000000000000000000111111;
mem_nr_5[28] <= 32'b00000000000000000000000000111111;
mem_nr_5[29] <= 32'b11111111111111111111111111111111;
mem_nr_5[30] <= 32'b11111111111111111111111111111111;
mem_nr_5[31] <= 32'b11111111111111111111111111111111;


mem_nr_6[0] <= 32'b11111111111111111111111111111111;
mem_nr_6[1] <= 32'b11111111111111111111111111111111;
mem_nr_6[2] <= 32'b11111111111111111111111111111111;
mem_nr_6[3] <= 32'b11111100000000000000000000000000;
mem_nr_6[4] <= 32'b11111100000000000000000000000000;
mem_nr_6[5] <= 32'b11111100000000000000000000000000;
mem_nr_6[6] <= 32'b11111100000000000000000000000000;
mem_nr_6[7] <= 32'b11111100000000000000000000000000;
mem_nr_6[8] <= 32'b11111100000000000000000000000000;
mem_nr_6[9] <= 32'b11111100000000000000000000000000;
mem_nr_6[10] <= 32'b11111100000000000000000000000000;
mem_nr_6[11] <= 32'b11111100000000000000000000000000;
mem_nr_6[12] <= 32'b11111100000000000000000000000000;
mem_nr_6[13] <= 32'b11111111111111111111111111111111;
mem_nr_6[14] <= 32'b11111111111111111111111111111111;
mem_nr_6[15] <= 32'b11111111111111111111111111111111;
mem_nr_6[16] <= 32'b11111111111111111111111111111111;
mem_nr_6[17] <= 32'b11111111111111111111111111111111;
mem_nr_6[18] <= 32'b11111100000000000000000000111111;
mem_nr_6[19] <= 32'b11111100000000000000000000111111;
mem_nr_6[20] <= 32'b11111100000000000000000000111111;
mem_nr_6[21] <= 32'b11111100000000000000000000111111;
mem_nr_6[22] <= 32'b11111100000000000000000000111111;
mem_nr_6[23] <= 32'b11111100000000000000000000111111;
mem_nr_6[24] <= 32'b11111100000000000000000000111111;
mem_nr_6[25] <= 32'b11111100000000000000000000111111;
mem_nr_6[26] <= 32'b11111100000000000000000000111111;
mem_nr_6[27] <= 32'b11111100000000000000000000111111;
mem_nr_6[28] <= 32'b11111100000000000000000000111111;
mem_nr_6[29] <= 32'b11111111111111111111111111111111;
mem_nr_6[30] <= 32'b11111111111111111111111111111111;
mem_nr_6[31] <= 32'b11111111111111111111111111111111;


mem_nr_7[0] <= 32'b11111111111111111111111111111111;
mem_nr_7[1] <= 32'b11111111111111111111111111111111;
mem_nr_7[2] <= 32'b11111111111111111111111111111111;
mem_nr_7[3] <= 32'b00000000000000000000000000111111;
mem_nr_7[4] <= 32'b00000000000000000000000000111111;
mem_nr_7[5] <= 32'b00000000000000000000000000111111;
mem_nr_7[6] <= 32'b00000000000000000000000000111111;
mem_nr_7[7] <= 32'b00000000000000000000000000111111;
mem_nr_7[8] <= 32'b00000000000000000000000000111111;
mem_nr_7[9] <= 32'b00000000000000000000000000111111;
mem_nr_7[10] <= 32'b00000000000000000000000000111111;
mem_nr_7[11] <= 32'b00000000000000000000000000111111;
mem_nr_7[12] <= 32'b00000000000000000000000000111111;
mem_nr_7[13] <= 32'b00000000000000000000000000111111;
mem_nr_7[14] <= 32'b00000000000000000000000000111111;
mem_nr_7[15] <= 32'b00000000000000000000000000111111;
mem_nr_7[16] <= 32'b00000000000000000000000000111111;
mem_nr_7[17] <= 32'b00000000000000000000000000111111;
mem_nr_7[18] <= 32'b00000000000000000000000000111111;
mem_nr_7[19] <= 32'b00000000000000000000000000111111;
mem_nr_7[20] <= 32'b00000000000000000000000000111111;
mem_nr_7[21] <= 32'b00000000000000000000000000111111;
mem_nr_7[22] <= 32'b00000000000000000000000000111111;
mem_nr_7[23] <= 32'b00000000000000000000000000111111;
mem_nr_7[24] <= 32'b00000000000000000000000000111111;
mem_nr_7[25] <= 32'b00000000000000000000000000111111;
mem_nr_7[26] <= 32'b00000000000000000000000000111111;
mem_nr_7[27] <= 32'b00000000000000000000000000111111;
mem_nr_7[28] <= 32'b00000000000000000000000000111111;
mem_nr_7[29] <= 32'b00000000000000000000000000111111;
mem_nr_7[30] <= 32'b00000000000000000000000000111111;
mem_nr_7[31] <= 32'b00000000000000000000000000111111;



mem_nr_8[0] <= 32'b11111111111111111111111111111111;
mem_nr_8[1] <= 32'b11111111111111111111111111111111;
mem_nr_8[2] <= 32'b11111111111111111111111111111111;
mem_nr_8[3] <= 32'b11111100000000000000000000111111;
mem_nr_8[4] <= 32'b11111100000000000000000000111111;
mem_nr_8[5] <= 32'b11111100000000000000000000111111;
mem_nr_8[6] <= 32'b11111100000000000000000000111111;
mem_nr_8[7] <= 32'b11111100000000000000000000111111;
mem_nr_8[8] <= 32'b11111100000000000000000000111111;
mem_nr_8[9] <= 32'b11111100000000000000000000111111;
mem_nr_8[10] <= 32'b11111100000000000000000000111111;
mem_nr_8[11] <= 32'b11111100000000000000000000111111;
mem_nr_8[12] <= 32'b11111100000000000000000000111111;
mem_nr_8[13] <= 32'b11111111111111111111111111111111;
mem_nr_8[14] <= 32'b11111111111111111111111111111111;
mem_nr_8[15] <= 32'b11111111111111111111111111111111;
mem_nr_8[16] <= 32'b11111111111111111111111111111111;
mem_nr_8[17] <= 32'b11111111111111111111111111111111;
mem_nr_8[18] <= 32'b11111100000000000000000000111111;
mem_nr_8[19] <= 32'b11111100000000000000000000111111;
mem_nr_8[20] <= 32'b11111100000000000000000000111111;
mem_nr_8[21] <= 32'b11111100000000000000000000111111;
mem_nr_8[22] <= 32'b11111100000000000000000000111111;
mem_nr_8[23] <= 32'b11111100000000000000000000111111;
mem_nr_8[24] <= 32'b11111100000000000000000000111111;
mem_nr_8[25] <= 32'b11111100000000000000000000111111;
mem_nr_8[26] <= 32'b11111100000000000000000000111111;
mem_nr_8[27] <= 32'b11111100000000000000000000111111;
mem_nr_8[28] <= 32'b11111100000000000000000000111111;
mem_nr_8[29] <= 32'b11111111111111111111111111111111;
mem_nr_8[30] <= 32'b11111111111111111111111111111111;
mem_nr_8[31] <= 32'b11111111111111111111111111111111;



mem_nr_9[0] <= 32'b11111111111111111111111111111111;
mem_nr_9[1] <= 32'b11111111111111111111111111111111;
mem_nr_9[2] <= 32'b11111111111111111111111111111111;
mem_nr_9[3] <= 32'b11111100000000000000000000111111;
mem_nr_9[4] <= 32'b11111100000000000000000000111111;
mem_nr_9[5] <= 32'b11111100000000000000000000111111;
mem_nr_9[6] <= 32'b11111100000000000000000000111111;
mem_nr_9[7] <= 32'b11111100000000000000000000111111;
mem_nr_9[8] <= 32'b11111100000000000000000000111111;
mem_nr_9[9] <= 32'b11111100000000000000000000111111;
mem_nr_9[10] <= 32'b11111100000000000000000000111111;
mem_nr_9[11] <= 32'b11111100000000000000000000111111;
mem_nr_9[12] <= 32'b11111100000000000000000000111111;
mem_nr_9[13] <= 32'b11111111111111111111111111111111;
mem_nr_9[14] <= 32'b11111111111111111111111111111111;
mem_nr_9[15] <= 32'b11111111111111111111111111111111;
mem_nr_9[16] <= 32'b11111111111111111111111111111111;
mem_nr_9[17] <= 32'b11111111111111111111111111111111;
mem_nr_9[18] <= 32'b00000000000000000000000000111111;
mem_nr_9[19] <= 32'b00000000000000000000000000111111;
mem_nr_9[20] <= 32'b00000000000000000000000000111111;
mem_nr_9[21] <= 32'b00000000000000000000000000111111;
mem_nr_9[22] <= 32'b00000000000000000000000000111111;
mem_nr_9[23] <= 32'b00000000000000000000000000111111;
mem_nr_9[24] <= 32'b00000000000000000000000000111111;
mem_nr_9[25] <= 32'b00000000000000000000000000111111;
mem_nr_9[26] <= 32'b00000000000000000000000000111111;
mem_nr_9[27] <= 32'b00000000000000000000000000111111;
mem_nr_9[28] <= 32'b00000000000000000000000000111111;
mem_nr_9[29] <= 32'b11111111111111111111111111111111;
mem_nr_9[30] <= 32'b11111111111111111111111111111111;
mem_nr_9[31] <= 32'b11111111111111111111111111111111;

    end
    else if(en_in) begin
        line_out_ff <= line_out_d;
    end
    else begin
        line_out_ff <= DISABLE;
    end
end

always @(*) begin
    line_out_d = line_out_ff;

    case (digit_in)

    ZERO: line_out_d = buffer_0;
    ONE: line_out_d = buffer_1;
    TWO: line_out_d = buffer_2;
    THREE: line_out_d = buffer_3;
    FOUR: line_out_d = buffer_4;
    FIVE: line_out_d = buffer_5;
    SIX: line_out_d = buffer_6;
    SEVEN: line_out_d = buffer_7;
    EIGTH: line_out_d = buffer_8;
    NINE: line_out_d = buffer_9;
        
        default: begin
            
        end
    endcase

end

assign line_out = line_out_ff;

assign buffer_0 = mem_nr_0[line_in];
assign buffer_1 = mem_nr_1[line_in];
assign buffer_2 = mem_nr_2[line_in];
assign buffer_3 = mem_nr_3[line_in];
assign buffer_4 = mem_nr_4[line_in];
assign buffer_5 = mem_nr_5[line_in];
assign buffer_6 = mem_nr_6[line_in];
assign buffer_7 = mem_nr_7[line_in];
assign buffer_8 = mem_nr_8[line_in];
assign buffer_9 = mem_nr_9[line_in];


endmodule