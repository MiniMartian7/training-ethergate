`include "sif_interface.sv"
`include "class_enviroment.sv"

module top;
    logic bit clk_top, rst_n_top;

    sif_interface top_i(clk_top);
    

endmodule : top