package lib_pack;
    typedef enum logic [2:0] {WRITE = 3'b110, READ = 3'b101, IDLE = 3'b100, ILLEGAL = 3'b111, RESET = 3'b000} E_Operation;
endpackage
/*aceasta este modificare ce trebuie sa apara in github*/
