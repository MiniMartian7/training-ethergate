module sif_tb;

sif_i tb_ports;
/*
modport TB (
        input clk,
        input xa_data_rd, wa_addr, wa_data_wr,
        output rst_n,
        output xa_addr, xa_data_wr,
        output xa_wr_s, xa_rd_s, wa_wr_s//enables
    );
*/




initial begin
    
end
endmodule