module mem(
    clk_mem,
    rst_mem,

    digit_in,

    pixel_out
);

input clk_mem, rst_mem;
input [3:0] digit_in;
output pixel_out;

reg [5:0] h_d, h_ff;
reg [5:0] v_d, v_ff;

reg pixel_buffer_d, pixel_buffer_ff;

reg display_block_d, display_block_ff;

reg [32:0] mem_nr_0 ;

reg [32:0] mem_nr_1 ;

reg [32:0] mem_nr_2; 

reg [32:0] mem_nr_3; 

reg [32:0] mem_nr_4; 

reg [32:0] mem_nr_5;

reg [32:0] mem_nr_6;

reg [32:0] mem_nr_7;

reg [32:0] mem_nr_8;

reg [32:0] mem_nr_9;

parameter ZERO = 'd0;
parameter ONE = 'd1;
parameter TWO = 'd2;
parameter THREE = 'd3;
parameter FOUR = 'd4;
parameter FIVE = 'd5;
parameter SIX = 'd6;
parameter SEVEN = 'd7;
parameter EIGTH = 'd8;
parameter NINE = 'd9;
parameter TEN = 'd10;

parameter NULL = 'b1111;

parameter ENABLE = 1;
parameter DISABLE = 0;
parameter RESET = 0;

always @(posedge clk_mem or posedge rst_mem) begin
    if(rst_mem) begin
        h_ff <= RESET;
        v_ff <=RESET;

        pixel_buffer_ff <= RESET; 

        display_block_ff <= RESET;     

        mem_nr_0 <= {
32'b11111111111111111111111111111111, 
32'b11111111111111111111111111111111, 
32'b11111111111111111111111111111111, 
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111111111111111111111111111111, 
32'b11111111111111111111111111111111, 
32'b11111111111111111111111111111111
};  

mem_nr_1 <= {
32'b00000000000000000000000111111111,
32'b00000000000000000000011111111111,
32'b00000000000000000001111111111111,
32'b00000000000000000111111111111111,
32'b00000000000000011111111100111111,
32'b00000000000001111111110000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111
};

mem_nr_2 <= {
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111
};

mem_nr_3 <= {
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111
};

mem_nr_4 <= {
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111
};

mem_nr_5 <= {
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111
};

mem_nr_6 <= {
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111
};

mem_nr_7 <= {
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111
};

mem_nr_8 <= {
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111
};

mem_nr_9 <= {
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111100000000000000000000111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b00000000000000000000000000111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111
};
    end
    else begin
        h_ff <= h_d;
        v_ff <= v_d;

        pixel_buffer_ff <= pixel_buffer_d;

        display_block_ff <= display_block_d;
    end
end

always @(*) begin
    h_d = h_ff;
    v_d = v_ff;

    pixel_buffer_d = pixel_buffer_ff;

    display_block_d = display_block_ff;

    if(display_block_ff == DISABLE) begin
        if(v_ff == 'd32) begin
            h_d = DISABLE;
            v_d = DISABLE;
            display_block_d = ENABLE;
        end
        else if(h_ff == 'd32) begin
            h_d = RESET;
            v_d = v_d + 1;
            display_block_d = ENABLE;
        end
        else begin
            h_d = h_d + 1;
        end
    end
    else begin
        h_d = DISABLE;
        v_d = DISABLE;
    end

    if(digit_in == ZERO) begin
        display_block_d = DISABLE;
        pixel_buffer_d = (mem_nr_0[v_d] << h_d ) & ('h80000000);
    end
    else if(digit_in == ONE) begin
        display_block_d = DISABLE;
        pixel_buffer_d = (mem_nr_1[v_d] << h_d ) & ('h80000000);
    end
    else if(digit_in == TWO) begin
        display_block_d = DISABLE;
        pixel_buffer_d = (mem_nr_2[v_d] << h_d ) & ('h80000000);
    end
    else if(digit_in == THREE) begin
        display_block_d = DISABLE;
        pixel_buffer_d = (mem_nr_3[v_d] << h_d ) & ('h80000000);
    end
    else if(digit_in == FOUR) begin
        display_block_d = DISABLE;
        pixel_buffer_d = (mem_nr_4[v_d] << h_d ) & ('h80000000);
    end
    else if(digit_in == FIVE) begin
        display_block_d = DISABLE;
        pixel_buffer_d = (mem_nr_5[v_d] << h_d ) & ('h80000000);
    end
    else if(digit_in == SIX) begin
        display_block_d = DISABLE;
        pixel_buffer_d = (mem_nr_6[v_d] << h_d ) & ('h80000000);
    end
    else if(digit_in == SEVEN) begin
        display_block_d = DISABLE;
        pixel_buffer_d = (mem_nr_7[v_d] << h_d ) & ('h80000000);
    end
    else if(digit_in == EIGTH) begin
        display_block_d = DISABLE;
        pixel_buffer_d = (mem_nr_8[v_d] << h_d ) & ('h80000000);
    end
    else if(digit_in == NINE) begin
        display_block_d = DISABLE;
        pixel_buffer_d = (mem_nr_9[v_d] << h_d ) & ('h80000000);
    end
    else if(digit_in == NULL) begin
        display_block_d = ENABLE;
        pixel_buffer_d = DISABLE;
    end
end

assign pixel_out = pixel_buffer_ff;

endmodule